`timescale 1ns / 1ps

module z1top(
  input a,
  input b,
  output c
);
  and(c, a, b);
endmodule
