`timescale 1ns/1ns

module structural_adder (
  input [2:0] a,
  input [2:0] b,
  output [3:0] sum
);
  // TODO: Insert your RTL here
  // Remove the assign statement once you write your own RTL
  assign sum = 4'd0;

endmodule
