
module uart #(
  parameter CLOCK_FREQ = 125_000_000,
  parameter BAUD_RATE  = 115_200
) (
  input clk,
  input rst,

  input  serial_in,
  output serial_out
);

  // TODO: Your code. Feel free to use any modules you like
  // Perform case inversion on letters only

endmodule
