`define BLACK   24'h000000
`define WHITE   24'hFFFFFF
`define GREEN   24'h00FF00
`define BLUE    24'h0000FF
`define RED     24'hFF0000
`define SILVER  24'hC0C0C0
`define GRAY    24'h808080
`define MAROON  24'h800000
`define YELLOW  24'hFFFF00
`define AQUA    24'h00FFFF
`define NAVY    24'h000080
`define MAGENTA 24'hFF00FF
`define TEAL    24'h008080
`define PURPLE  24'h800080
